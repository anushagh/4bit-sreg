//transactor class

class transactor;

rand bit serial_in;
rand bit [3:0] parallel_in;
rand bit dir,load;

endclass
